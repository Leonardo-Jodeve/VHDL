-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 9.0 Build 132 02/25/2009 SJ Full Version"
-- CREATED ON		"Mon Sep 07 22:29:28 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY TrafficLight IS 
	PORT
	(
		pin_name :  IN  STD_LOGIC;
		Main_Red :  OUT  STD_LOGIC;
		Main_Yellow :  OUT  STD_LOGIC;
		Main_Green :  OUT  STD_LOGIC;
		Vice_Red :  OUT  STD_LOGIC;
		Vice_Yellow :  OUT  STD_LOGIC;
		Vice_Green :  OUT  STD_LOGIC
	);
END TrafficLight;

ARCHITECTURE bdf_type OF TrafficLight IS 

ATTRIBUTE black_box : BOOLEAN;
nATTRIBUTE noopt : BOOLEAN;

COMPONENT \74160_0\
	PORT(CLK : IN STD_LOGIC;
		 ENT : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 LDN : IN STD_LOGIC;
		 ENP : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74160_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \74160_0\: COMPONENT IS true;

COMPONENT \74190_1\
	PORT(A : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 RCON : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74190_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \74190_1\: COMPONENT IS true;

COMPONENT \74190_2\
	PORT(A : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 MXMN : OUT STD_LOGIC;
		 RCON : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74190_2\: COMPONENT IS true;
ATTRIBUTE noopt OF \74190_2\: COMPONENT IS true;

COMPONENT \74190_3\
	PORT(A : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 RCON : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74190_3\: COMPONENT IS true;
ATTRIBUTE noopt OF \74190_3\: COMPONENT IS true;

COMPONENT \74190_4\
	PORT(A : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 DNUP : IN STD_LOGIC;
		 MXMN : OUT STD_LOGIC;
		 RCON : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74190_4\: COMPONENT IS true;
ATTRIBUTE noopt OF \74190_4\: COMPONENT IS true;

SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;


BEGIN 
Main_Yellow <= SYNTHESIZED_WIRE_55;
Main_Green <= SYNTHESIZED_WIRE_56;
Vice_Yellow <= SYNTHESIZED_WIRE_49;
Vice_Green <= SYNTHESIZED_WIRE_50;
SYNTHESIZED_WIRE_53 <= '1';
SYNTHESIZED_WIRE_54 <= '0';
SYNTHESIZED_WIRE_57 <= '0';
SYNTHESIZED_WIRE_59 <= '0';



SYNTHESIZED_WIRE_60 <= SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_50;


SYNTHESIZED_WIRE_56 <= NOT(SYNTHESIZED_WIRE_51 OR SYNTHESIZED_WIRE_52);


SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_4 AND SYNTHESIZED_WIRE_51;


SYNTHESIZED_WIRE_4 <= NOT(SYNTHESIZED_WIRE_52);



SYNTHESIZED_WIRE_50 <= SYNTHESIZED_WIRE_52 AND SYNTHESIZED_WIRE_8;


SYNTHESIZED_WIRE_8 <= NOT(SYNTHESIZED_WIRE_51);



SYNTHESIZED_WIRE_49 <= SYNTHESIZED_WIRE_52 AND SYNTHESIZED_WIRE_51;



b2v_inst21 : 74160_0
PORT MAP(CLK => SYNTHESIZED_WIRE_12,
		 ENT => SYNTHESIZED_WIRE_53,
		 A => SYNTHESIZED_WIRE_54,
		 B => SYNTHESIZED_WIRE_54,
		 C => SYNTHESIZED_WIRE_54,
		 D => SYNTHESIZED_WIRE_54,
		 LDN => SYNTHESIZED_WIRE_18,
		 ENP => SYNTHESIZED_WIRE_53,
		 CLRN => SYNTHESIZED_WIRE_53,
		 QA => SYNTHESIZED_WIRE_52,
		 QB => SYNTHESIZED_WIRE_51,
		 QC => SYNTHESIZED_WIRE_18);



Main_Red <= SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_50;


Vice_Red <= SYNTHESIZED_WIRE_55 OR SYNTHESIZED_WIRE_56;


b2v_inst34 : 74190_1
PORT MAP(A => SYNTHESIZED_WIRE_50,
		 C => SYNTHESIZED_WIRE_56,
		 B => SYNTHESIZED_WIRE_50,
		 CLK => SYNTHESIZED_WIRE_28,
		 DNUP => SYNTHESIZED_WIRE_57,
		 RCON => SYNTHESIZED_WIRE_41);


b2v_inst35 : 74190_2
PORT MAP(A => SYNTHESIZED_WIRE_58,
		 C => SYNTHESIZED_WIRE_58,
		 CLK => pin_name,
		 DNUP => SYNTHESIZED_WIRE_57,
		 MXMN => SYNTHESIZED_WIRE_28,
		 RCON => SYNTHESIZED_WIRE_42);


b2v_inst36 : 74190_3
PORT MAP(A => SYNTHESIZED_WIRE_56,
		 C => SYNTHESIZED_WIRE_56,
		 B => SYNTHESIZED_WIRE_50,
		 CLK => SYNTHESIZED_WIRE_36,
		 DNUP => SYNTHESIZED_WIRE_59,
		 RCON => SYNTHESIZED_WIRE_43);


b2v_inst37 : 74190_4
PORT MAP(A => SYNTHESIZED_WIRE_60,
		 C => SYNTHESIZED_WIRE_60,
		 CLK => pin_name,
		 DNUP => SYNTHESIZED_WIRE_59,
		 MXMN => SYNTHESIZED_WIRE_36,
		 RCON => SYNTHESIZED_WIRE_44);




SYNTHESIZED_WIRE_47 <= SYNTHESIZED_WIRE_41 OR SYNTHESIZED_WIRE_42;


SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_43 OR SYNTHESIZED_WIRE_44;


SYNTHESIZED_WIRE_58 <= SYNTHESIZED_WIRE_56 OR SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_47 OR SYNTHESIZED_WIRE_48;


END bdf_type;